* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_76_199# a_206_369# a_489_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR a_206_369# a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 VPWR A1_N a_206_369# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_206_369# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VGND B1 a_489_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 X a_76_199# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_489_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 X a_76_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X8 a_205_47# A2_N a_206_369# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_76_199# B2 a_585_369# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_585_369# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 VGND A1_N a_205_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
