* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
X0 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X1 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X3 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X4 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X5 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X6 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X7 a_465_47# B a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_27_47# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X10 a_215_47# B a_465_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_655_47# C a_465_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VGND D a_655_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_27_47# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_465_47# C a_655_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_655_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
.ends
