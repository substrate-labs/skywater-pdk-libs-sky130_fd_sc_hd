* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 a_136_47# B2 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VPWR B2 a_54_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X2 a_442_21# A2_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 Y a_442_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VGND A2_N a_442_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VGND A1_N a_442_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_54_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X7 VGND a_442_21# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_662_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X9 a_442_21# A1_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_136_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VPWR B1 a_54_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X12 VPWR A1_N a_662_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X13 Y a_442_21# a_54_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X14 a_442_21# A2_N a_662_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X15 Y B2 a_136_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_54_297# B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X17 VGND B1 a_136_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_54_297# a_442_21# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X19 a_662_297# A2_N a_442_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
.ends
