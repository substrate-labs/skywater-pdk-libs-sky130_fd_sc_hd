* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
X0 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_542_297# B a_626_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_626_297# a_27_47# a_176_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X5 a_27_47# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND A a_176_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X9 a_27_47# C_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X11 VGND a_27_47# a_176_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X13 VPWR A a_542_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X14 a_176_21# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
.ends
