* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_4 A LOWLVPWR VGND VNB VPB VPWR X
X0 a_424_82# a_1032_911# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 X a_1032_911# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X2 VPWR a_1032_911# X VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X3 X a_1032_911# a_424_82# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_714_47# a_620_911# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X5 a_620_911# a_505_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_620_911# a_505_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 X a_1032_911# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X8 a_424_82# A a_714_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 LOWLVPWR A a_505_297# LOWLVPWR sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X10 a_714_47# A a_424_82# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VPWR a_1032_911# X VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X12 VPWR a_620_911# a_1032_911# VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X13 a_424_82# a_1032_911# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VGND a_505_297# a_620_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 X a_1032_911# a_424_82# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VGND a_505_297# a_620_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_424_82# A a_714_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_714_47# A a_424_82# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 VGND a_620_911# a_1032_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_620_911# a_714_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=790000u l=150000u
X21 a_424_82# A a_505_297# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
