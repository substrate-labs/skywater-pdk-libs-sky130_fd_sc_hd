* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
X0 VPWR A1 a_1243_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X1 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VGND A4 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VGND A4 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_467_297# A4 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X7 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 Y A4 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X10 a_885_297# A2 a_1243_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X11 a_885_297# A2 a_1243_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X12 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_885_297# A3 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X15 VPWR A1 a_1243_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X16 a_1243_297# A2 a_885_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X17 a_27_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_467_297# A3 a_885_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X19 a_1243_297# A2 a_885_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X20 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_27_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 a_1243_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X25 a_885_297# A3 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X26 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X29 a_467_297# A4 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X30 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 a_467_297# A3 a_885_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X32 a_1243_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X33 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X34 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X35 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X36 Y A4 a_467_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X37 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X38 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X39 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
