* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__nand4bb_1 A_N B_N C D VGND VNB VPB VPWR Y
X0 Y a_496_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X1 a_426_47# a_496_21# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR A_N a_496_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 VGND A_N a_496_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_27_93# B_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X6 a_326_47# a_27_93# a_426_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_27_93# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X9 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X10 VGND D a_218_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_218_47# C a_326_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
