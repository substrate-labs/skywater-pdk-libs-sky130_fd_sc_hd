* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
X0 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X3 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_193_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X8 a_27_47# C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_27_47# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X11 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X12 a_109_297# B a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1 l=150000u
X13 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
